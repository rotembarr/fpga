package multiply_pack;
	typedef enum int {
		DSP,
		LUTS
	} multiply_t;

	typedef enum int {
		LOGIC,
		LUTS
	} signed_add_t;
endpackage